`timescale 1ns / 1ps


module SPI_test;

	// Outputs
	wire ;

	// Instantiate the Unit Under Test (UUT)
	SPI_Master uut (
		.()
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here

	end
      
endmodule

